module test_simple (input logic clk); logic [7:0] test; endmodule
